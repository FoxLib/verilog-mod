`timescale 10ns / 1ns
module tb;
// ---------------------------------------------------------------------
reg clock;
reg clock_25;
reg clock_50;

always #0.5 clock    = ~clock;
always #1.0 clock_50 = ~clock_50;
always #1.5 clock_25 = ~clock_25;

initial begin clock = 1; clock_25 = 0; clock_50 = 0; #2000 $finish; end
initial begin $dumpfile("tb.vcd"); $dumpvars(0, tb); end
// ---------------------------------------------------------------------

wire cs;
wire sclk;
wire miso;
wire mosi;

sdcard SD(

    .clock      (clock),
    .spi_cs     (cs),
    .spi_sclk   (sclk),
    .spi_miso   (miso),
    .spi_mosi   (mosi)
);

endmodule
